module Flags(
    input [2:0] alu_iFlags,
    output [2:0] oFlags_uc
    );
endmodule